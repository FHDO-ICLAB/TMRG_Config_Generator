
class rdc;
    int rdc_success ,rdc_fail;

    function new;
        this.rdc_success = $fopen("./rdc_success.txt", "w");
        this.rdc_fail = $fopen("./rdc_fail.txt", "w");
    endfunction

    function logging(string func,string add, string msg);
        if (func == add) begin
            $fdisplay(this.rdc_success, "%s", msg);
        end else begin
            $fdisplay(this.rdc_success, "%s", msg);
        end
    endfunction
    
    function reset(string appendix);
        case (appendix)
            "A" : this.resetA;
            "B" : this.resetB;
            "C" : this.resetC;
            default : $stop;
        endcase
    endfunction
    
    function resetA;
        assert(top_test.can2TMR_u.TimeControl.smpldbit_reg_i.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.smpldbit_reg_i.resetA");

		assert(top_test.can2TMR_u.TimeControl.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.resetA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.pid_regler0.OutputScaling0.ResetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.pid_regler0.OutputScaling0.ResetA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.control_fsm0.ResetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.control_fsm0.ResetA");

		assert(top_test.can2TMR_u.TimeControl.bittiming.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.bittiming.resetA");

		assert(top_test.can2TMR_u.reset_generator.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.reset_generator.resetA");

		assert(top_test.can2TMR_u.prescaler.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.prescaler.resetA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[14].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[14].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[13].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[13].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[12].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[12].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[11].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[11].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[10].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[10].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[9].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[9].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[8].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[8].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[7].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[7].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[6].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[6].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[5].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[5].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[4].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[4].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[3].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[3].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[2].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[2].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[1].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[1].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[0].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[0].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.activ_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.activ_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.topreg.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.topreg.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[101].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[101].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[100].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[100].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[99].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[99].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[98].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[98].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[97].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[97].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[96].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[96].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[95].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[95].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[94].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[94].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[93].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[93].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[92].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[92].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[91].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[91].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[90].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[90].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[89].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[89].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[88].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[88].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[87].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[87].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[86].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[86].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[85].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[85].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[84].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[84].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[83].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[83].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[82].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[82].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[81].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[81].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[80].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[80].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[79].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[79].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[78].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[78].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[77].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[77].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[76].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[76].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[75].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[75].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[74].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[74].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[73].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[73].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[72].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[72].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[71].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[71].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[70].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[70].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[69].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[69].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[68].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[68].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[67].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[67].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[66].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[66].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[65].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[65].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[64].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[64].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[63].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[63].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[62].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[62].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[61].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[61].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[60].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[60].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[59].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[59].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[58].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[58].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[57].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[57].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[56].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[56].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[55].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[55].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[54].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[54].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[53].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[53].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[52].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[52].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[51].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[51].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[50].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[50].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[49].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[49].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[48].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[48].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[47].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[47].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[46].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[46].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[45].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[45].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[44].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[44].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[43].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[43].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[42].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[42].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[41].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[41].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[40].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[40].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[39].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[39].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[38].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[38].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[37].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[37].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[36].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[36].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[35].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[35].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[34].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[34].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[33].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[33].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[32].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[32].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[31].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[31].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[30].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[30].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[29].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[29].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[28].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[28].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[27].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[27].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[26].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[26].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[25].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[25].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[24].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[24].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[23].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[23].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[22].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[22].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[21].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[21].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[20].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[20].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[19].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[19].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[18].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[18].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[17].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[17].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[16].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[16].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[15].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[15].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[14].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[14].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[13].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[13].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[12].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[12].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[11].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[11].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[10].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[10].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[9].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[9].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[8].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[8].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[7].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[7].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[6].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[6].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[5].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[5].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[4].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[4].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[3].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[3].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[2].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[2].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[1].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[1].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.enable_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.enable_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.bottom_reg.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.bottom_reg.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.stuff_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.stuff_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.BufA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.BufA");

		assert(top_test.can2TMR_u.MediumAccessControl.reset_mac_i.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.reset_mac_i.resetA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[102].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[102].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[101].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[101].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[100].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[100].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[99].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[99].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[98].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[98].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[97].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[97].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[96].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[96].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[95].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[95].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[94].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[94].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[93].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[93].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[92].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[92].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[91].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[91].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[90].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[90].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[89].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[89].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[88].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[88].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[87].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[87].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[86].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[86].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[85].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[85].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[84].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[84].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[83].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[83].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[82].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[82].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[81].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[81].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[80].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[80].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[79].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[79].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[78].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[78].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[77].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[77].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[76].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[76].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[75].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[75].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[74].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[74].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[73].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[73].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[72].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[72].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[71].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[71].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[70].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[70].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[69].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[69].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[68].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[68].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[67].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[67].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[66].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[66].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[65].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[65].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[64].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[64].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[63].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[63].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[62].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[62].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[61].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[61].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[60].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[60].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[59].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[59].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[58].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[58].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[57].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[57].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[56].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[56].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[55].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[55].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[54].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[54].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[53].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[53].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[52].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[52].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[51].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[51].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[50].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[50].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[49].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[49].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[48].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[48].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[47].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[47].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[46].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[46].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[45].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[45].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[44].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[44].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[43].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[43].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[42].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[42].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[41].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[41].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[40].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[40].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[39].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[39].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[38].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[38].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[37].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[37].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[36].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[36].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[35].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[35].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[34].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[34].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[33].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[33].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[32].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[32].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[31].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[31].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[30].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[30].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[29].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[29].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[28].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[28].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[27].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[27].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[26].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[26].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[25].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[25].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[24].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[24].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[23].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[23].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[22].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[22].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[21].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[21].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[20].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[20].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[19].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[19].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[18].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[18].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[17].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[17].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[16].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[16].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[15].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[15].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[14].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[14].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[13].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[13].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[12].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[12].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[11].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[11].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[10].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[10].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[9].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[9].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[8].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[8].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[7].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[7].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[6].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[6].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[5].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[5].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[4].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[4].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[3].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[3].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[2].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[2].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[1].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[1].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.enable_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.enable_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.bottom.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.bottom.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recmlen.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recmlen.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.transmitter_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.transmitter_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.rrtr_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.rrtr_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.rext_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.rext_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.receiver_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.receiver_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.puffer_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.puffer_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.first_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.first_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.error_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.error_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.ackerror_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.ackerror_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.workingA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.workingA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.directshift_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.directshift_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.errordetect.errorA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.errordetect.errorA");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.remA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.remA");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stuff_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stuff_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stfer_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stfer_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.inc_rise_merkerA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.inc_rise_merkerA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA");

		assert(top_test.can2TMR_u.irqunit.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.irqunit.CURRENT_STATEA");

		assert(top_test.can2TMR_u.irqunit.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.irqunit.CURRENT_STATEA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.edgedA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.edgedA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA");

		assert(top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA");

		assert(top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.edgedA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");
    endfunction

    function resetB;
        assert(top_test.can2TMR_u.TimeControl.smpldbit_reg_i.resetB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.smpldbit_reg_i.resetB");

		assert(top_test.can2TMR_u.TimeControl.resetB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.resetB");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnB");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnB");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnB");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnB");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnB");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.pid_regler0.OutputScaling0.ResetB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.pid_regler0.OutputScaling0.ResetB");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.control_fsm0.ResetB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.control_fsm0.ResetB");

		assert(top_test.can2TMR_u.TimeControl.bittiming.resetB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.bittiming.resetB");

		assert(top_test.can2TMR_u.reset_generator.resetB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.reset_generator.resetB");

		assert(top_test.can2TMR_u.prescaler.resetB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.prescaler.resetB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[14].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[14].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[13].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[13].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[12].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[12].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[11].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[11].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[10].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[10].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[9].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[9].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[8].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[8].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[7].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[7].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[6].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[6].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[5].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[5].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[4].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[4].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[3].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[3].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[2].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[2].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[1].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[1].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[0].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[0].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.activ_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.activ_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.edgedB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.edgedB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.topreg.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.topreg.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[101].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[101].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[100].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[100].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[99].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[99].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[98].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[98].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[97].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[97].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[96].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[96].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[95].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[95].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[94].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[94].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[93].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[93].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[92].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[92].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[91].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[91].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[90].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[90].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[89].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[89].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[88].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[88].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[87].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[87].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[86].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[86].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[85].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[85].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[84].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[84].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[83].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[83].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[82].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[82].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[81].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[81].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[80].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[80].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[79].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[79].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[78].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[78].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[77].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[77].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[76].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[76].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[75].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[75].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[74].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[74].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[73].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[73].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[72].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[72].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[71].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[71].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[70].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[70].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[69].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[69].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[68].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[68].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[67].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[67].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[66].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[66].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[65].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[65].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[64].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[64].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[63].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[63].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[62].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[62].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[61].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[61].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[60].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[60].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[59].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[59].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[58].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[58].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[57].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[57].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[56].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[56].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[55].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[55].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[54].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[54].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[53].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[53].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[52].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[52].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[51].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[51].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[50].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[50].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[49].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[49].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[48].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[48].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[47].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[47].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[46].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[46].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[45].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[45].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[44].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[44].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[43].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[43].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[42].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[42].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[41].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[41].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[40].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[40].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[39].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[39].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[38].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[38].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[37].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[37].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[36].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[36].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[35].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[35].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[34].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[34].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[33].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[33].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[32].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[32].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[31].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[31].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[30].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[30].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[29].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[29].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[28].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[28].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[27].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[27].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[26].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[26].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[25].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[25].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[24].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[24].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[23].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[23].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[22].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[22].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[21].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[21].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[20].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[20].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[19].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[19].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[18].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[18].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[17].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[17].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[16].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[16].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[15].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[15].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[14].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[14].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[13].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[13].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[12].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[12].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[11].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[11].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[10].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[10].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[9].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[9].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[8].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[8].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[7].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[7].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[6].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[6].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[5].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[5].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[4].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[4].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[3].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[3].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[2].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[2].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[1].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[1].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.enable_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.enable_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.edgedB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.edgedB");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.bottom_reg.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.bottom_reg.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.stuff_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.stuff_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.edgedB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.edgedB");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.BufB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.BufB");

		assert(top_test.can2TMR_u.MediumAccessControl.reset_mac_i.resetB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.reset_mac_i.resetB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[102].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[102].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[101].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[101].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[100].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[100].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[99].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[99].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[98].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[98].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[97].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[97].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[96].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[96].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[95].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[95].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[94].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[94].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[93].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[93].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[92].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[92].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[91].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[91].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[90].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[90].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[89].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[89].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[88].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[88].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[87].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[87].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[86].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[86].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[85].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[85].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[84].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[84].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[83].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[83].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[82].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[82].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[81].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[81].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[80].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[80].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[79].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[79].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[78].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[78].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[77].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[77].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[76].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[76].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[75].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[75].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[74].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[74].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[73].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[73].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[72].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[72].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[71].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[71].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[70].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[70].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[69].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[69].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[68].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[68].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[67].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[67].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[66].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[66].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[65].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[65].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[64].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[64].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[63].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[63].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[62].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[62].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[61].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[61].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[60].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[60].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[59].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[59].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[58].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[58].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[57].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[57].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[56].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[56].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[55].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[55].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[54].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[54].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[53].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[53].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[52].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[52].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[51].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[51].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[50].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[50].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[49].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[49].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[48].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[48].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[47].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[47].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[46].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[46].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[45].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[45].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[44].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[44].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[43].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[43].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[42].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[42].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[41].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[41].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[40].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[40].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[39].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[39].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[38].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[38].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[37].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[37].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[36].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[36].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[35].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[35].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[34].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[34].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[33].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[33].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[32].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[32].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[31].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[31].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[30].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[30].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[29].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[29].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[28].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[28].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[27].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[27].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[26].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[26].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[25].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[25].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[24].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[24].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[23].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[23].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[22].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[22].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[21].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[21].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[20].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[20].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[19].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[19].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[18].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[18].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[17].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[17].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[16].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[16].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[15].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[15].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[14].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[14].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[13].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[13].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[12].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[12].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[11].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[11].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[10].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[10].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[9].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[9].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[8].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[8].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[7].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[7].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[6].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[6].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[5].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[5].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[4].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[4].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[3].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[3].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[2].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[2].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[1].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[1].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.enable_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.enable_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.edgedB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.edgedB");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.bottom.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.bottom.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.recmlen.edgedB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recmlen.edgedB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.q_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.q_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.edge_varB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.edge_varB");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.transmitter_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.transmitter_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.rrtr_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.rrtr_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.rext_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.rext_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.receiver_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.receiver_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.puffer_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.puffer_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.first_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.first_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.error_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.error_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.ackerror_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.ackerror_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.workingB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.workingB");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.directshift_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.directshift_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.errordetect.errorB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.errordetect.errorB");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.remB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.remB");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufB");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufB");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufB");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufB");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stuff_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stuff_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stfer_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stfer_iB");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateB");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateB");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateB");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateB");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.edgedB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.edgedB");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.inc_rise_merkerB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.inc_rise_merkerB");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countB");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countB");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEB");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEB");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEB");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEB");

		assert(top_test.can2TMR_u.irqunit.CURRENT_STATEB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.irqunit.CURRENT_STATEB");

		assert(top_test.can2TMR_u.irqunit.CURRENT_STATEB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.irqunit.CURRENT_STATEB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.general.register_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iB");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.edgedB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.edgedB");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.edgedB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.edgedB");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEB");

		assert(top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEB");

		assert(top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEB");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.edgedB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.edgedB");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterB");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterB)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterB");
    endfunction

    function resetC;
        assert(top_test.can2TMR_u.TimeControl.smpldbit_reg_i.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.smpldbit_reg_i.resetA");

		assert(top_test.can2TMR_u.TimeControl.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.resetA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.rdy_cnt0.rstnA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.pid_regler0.OutputScaling0.ResetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.pid_regler0.OutputScaling0.ResetA");

		assert(top_test.can2TMR_u.TimeControl.freqTrim.control_fsm0.ResetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.freqTrim.control_fsm0.ResetA");

		assert(top_test.can2TMR_u.TimeControl.bittiming.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.TimeControl.bittiming.resetA");

		assert(top_test.can2TMR_u.reset_generator.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.reset_generator.resetA");

		assert(top_test.can2TMR_u.prescaler.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.prescaler.resetA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[14].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[14].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[13].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[13].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[12].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[12].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[11].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[11].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[10].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[10].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[9].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[9].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[8].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[8].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[7].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[7].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[6].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[6].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[5].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[5].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[4].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[4].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[3].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[3].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[2].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[2].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[1].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[1].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[0].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.genblk1[0].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.activ_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.activ_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transmitcrc.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transmitcrc.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.topreg.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.topreg.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[101].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[101].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[100].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[100].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[99].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[99].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[98].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[98].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[97].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[97].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[96].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[96].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[95].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[95].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[94].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[94].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[93].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[93].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[92].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[92].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[91].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[91].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[90].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[90].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[89].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[89].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[88].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[88].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[87].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[87].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[86].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[86].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[85].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[85].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[84].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[84].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[83].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[83].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[82].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[82].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[81].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[81].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[80].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[80].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[79].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[79].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[78].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[78].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[77].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[77].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[76].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[76].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[75].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[75].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[74].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[74].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[73].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[73].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[72].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[72].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[71].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[71].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[70].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[70].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[69].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[69].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[68].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[68].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[67].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[67].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[66].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[66].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[65].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[65].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[64].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[64].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[63].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[63].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[62].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[62].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[61].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[61].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[60].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[60].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[59].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[59].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[58].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[58].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[57].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[57].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[56].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[56].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[55].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[55].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[54].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[54].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[53].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[53].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[52].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[52].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[51].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[51].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[50].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[50].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[49].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[49].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[48].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[48].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[47].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[47].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[46].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[46].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[45].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[45].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[44].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[44].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[43].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[43].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[42].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[42].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[41].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[41].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[40].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[40].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[39].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[39].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[38].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[38].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[37].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[37].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[36].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[36].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[35].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[35].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[34].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[34].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[33].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[33].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[32].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[32].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[31].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[31].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[30].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[30].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[29].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[29].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[28].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[28].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[27].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[27].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[26].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[26].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[25].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[25].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[24].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[24].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[23].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[23].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[22].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[22].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[21].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[21].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[20].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[20].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[19].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[19].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[18].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[18].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[17].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[17].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[16].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[16].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[15].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[15].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[14].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[14].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[13].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[13].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[12].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[12].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[11].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[11].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[10].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[10].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[9].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[9].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[8].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[8].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[7].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[7].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[6].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[6].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[5].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[5].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[4].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[4].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[3].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[3].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[2].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[2].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[1].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.genblk1[1].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.enable_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.enable_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.transhift.bottom_reg.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.transhift.bottom_reg.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.stuff_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.stuff_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.stuff.BufA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.stuff.BufA");

		assert(top_test.can2TMR_u.MediumAccessControl.reset_mac_i.resetA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.reset_mac_i.resetA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[102].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[102].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[101].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[101].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[100].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[100].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[99].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[99].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[98].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[98].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[97].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[97].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[96].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[96].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[95].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[95].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[94].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[94].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[93].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[93].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[92].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[92].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[91].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[91].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[90].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[90].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[89].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[89].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[88].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[88].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[87].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[87].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[86].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[86].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[85].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[85].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[84].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[84].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[83].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[83].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[82].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[82].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[81].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[81].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[80].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[80].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[79].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[79].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[78].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[78].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[77].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[77].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[76].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[76].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[75].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[75].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[74].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[74].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[73].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[73].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[72].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[72].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[71].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[71].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[70].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[70].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[69].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[69].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[68].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[68].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[67].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[67].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[66].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[66].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[65].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[65].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[64].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[64].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[63].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[63].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[62].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[62].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[61].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[61].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[60].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[60].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[59].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[59].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[58].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[58].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[57].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[57].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[56].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[56].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[55].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[55].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[54].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[54].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[53].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[53].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[52].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[52].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[51].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[51].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[50].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[50].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[49].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[49].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[48].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[48].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[47].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[47].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[46].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[46].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[45].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[45].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[44].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[44].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[43].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[43].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[42].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[42].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[41].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[41].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[40].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[40].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[39].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[39].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[38].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[38].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[37].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[37].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[36].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[36].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[35].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[35].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[34].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[34].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[33].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[33].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[32].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[32].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[31].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[31].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[30].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[30].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[29].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[29].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[28].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[28].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[27].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[27].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[26].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[26].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[25].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[25].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[24].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[24].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[23].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[23].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[22].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[22].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[21].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[21].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[20].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[20].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[19].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[19].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[18].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[18].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[17].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[17].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[16].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[16].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[15].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[15].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[14].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[14].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[13].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[13].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[12].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[12].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[11].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[11].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[10].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[10].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[9].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[9].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[8].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[8].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[7].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[7].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[6].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[6].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[5].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[5].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[4].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[4].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[3].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[3].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[2].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[2].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[1].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.genblk1[1].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.enable_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.enable_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.recshift.bottom.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recshift.bottom.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.recmlen.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.recmlen.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[14].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[13].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[12].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[11].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[10].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[9].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[8].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[7].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[6].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[5].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[4].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[3].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[2].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[1].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.q_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.q_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.edge_varA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.receivecrc.genblk1[0].reg_i.edge_varA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.transmitter_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.transmitter_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.rrtr_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.rrtr_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.rext_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.rext_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.receiver_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.receiver_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.puffer_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.puffer_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.first_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.first_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.error_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.error_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.fsm_regs.ackerror_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.fsm_regs.ackerror_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.workingA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.workingA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.directshift_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.directshift_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.frshift.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.frshift.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.errordetect.errorA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.errordetect.errorA");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.remA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.remA");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA");

		assert(top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.encaps.datalen_bufA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stuff_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stuff_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stfer_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stfer_iA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.stateA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.stateA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.edgedA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.destuff.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.destuff.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.inc_rise_merkerA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.inc_rise_merkerA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.MediumAccessControl.counting.countA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.MediumAccessControl.counting.countA");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA");

		assert(top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.LogicalLinkControl.llc_fsm_2.CURRENT_STATEA");

		assert(top_test.can2TMR_u.irqunit.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.irqunit.CURRENT_STATEA");

		assert(top_test.can2TMR_u.irqunit.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.irqunit.CURRENT_STATEA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.tarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.tarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata78.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata78.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata56.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata56.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata34.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata34.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rdata12.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rdata12.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit2.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit2.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.rarbit1.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.rarbit1.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.prescaleregister.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.prescaleregister.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.mcontrol.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.mcontrol.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.interruptreg.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.interruptreg.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.general.register_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.general.register_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask2.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask2.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.IOControl.accmask1.reg_iA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.IOControl.accmask1.reg_iA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.edgedA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.tec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.tec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.edgedA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.rec_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.rec_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA");

		assert(top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA");

		assert(top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.fsm.CURRENT_STATEA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.edgedA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.edgedA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");

		assert(top_test.can2TMR_u.FaultConfinement.erb_count.counterA)
		else
			$fdisplay(this.rdc_fail, "top_test.can2TMR_u.FaultConfinement.erb_count.counterA");
    endfunction
endclass    
